module bindfiles;
	bind lc3 lc3_asserts p1 (.*);
endmodule
