module bindfiles;
	bind lc3 lc3_asserts p1 (.*);
	bind regfile8x16 regfile_asserts p2 (.*);
endmodule
