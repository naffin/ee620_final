module bindfiles;
	bind top lc3_asserts p1 (.*);
endmodule
