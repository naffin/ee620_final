package svm_component_pkg;
virtual class svm_component;
	pure virtual task run_test();
endclass // svm_component_pkg
endpackage
