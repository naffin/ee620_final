package Coverage_base_pkg;
   import Transaction_pkg::*;
virtual class Coverage_base;
   pure virtual function void sample(Transaction t);
endclass
endpackage
   
