module bindfiles;
   bind datapath datapath_asserts dp_a(.*);
   bind controller controller_asserts fsm_a(.*);
endmodule
